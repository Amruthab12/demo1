//simple class example

class a;
	int [31:00] addr;
	bit id;

	function void display();
        $display("class example");
endfunction
endclass

